library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity p_enemy is
    port(
        x_e,y_e: in std_logic_vector(5 downto 0); --the xy for the plane and the enemy 
        d_e: out std_logic 
    );
end p_enemy;

architecture Behav of p_enemy is
    type d_block is array(0 to 31) of std_logic_vector(31 downto 0);
constant e_block: d_block :=
    ("11111111111111111111111111111111",
     "11111111111111111111111111111111",
     "11111111111111111111111111111111",
     "11111111111111111111111111111111",
     "11111111111111111111111111111111",
     "11111111111111111111111111111111",
     "11111111111111111111111111111111",
     "11111011111111111111111111011111",
     "11111011111111111111111111011111",
     "11111011111111111111111111011111",
     "11111011111111111111111111011111",
     "00000000000000000000000000000000",
     "00000000000000000000000000000000",
     "00000000000000000000000000000000",
     "01100000000000000000000000000110",
     "01111100000000000000000001111110",
     "01111111100000000000000111111110",
     "11111111111100000000111111111111",
     "11111111111110000001111111111111",
     "11111111111110000001111111111111",
     "11111111111111000011111111111111",
     "11111111111111000011111111111111",
     "11111111111111100111111111111111",
     "11111111111111100111111111111111",
     "11111111111111111111111111111111",
     "11111111111111111111111111111111",
     "11111111111111111111111111111111",
     "11111111111111111111111111111111",
     "11111111111111111111111111111111",
     "11111111111111111111111111111111",
     "11111111111111111111111111111111", 
     "11111111111111111111111111111111" );


signal tmp_e:std_logic_vector(31 downto 0);
begin 
tmp_e<=e_block(conv_integer(y_e));
d_e<=not tmp_e(conv_integer(x_e));
end Behav;